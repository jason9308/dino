module dino_crtl(
    input	lcd_pclk,
    input	rst_n,
    input	[10:0]  pixel_xpos,
    input	[10:0]  pixel_ypos, 
	input	key_flag,
	input	key_value,
	input	is_living,
	input	is_dying,
	
    output	dino_draw,
	output reg clk_100
);

/* --------------------------------------------------------------------------------------------------------------------------- */
	 
	reg [82:0] body_normal [73:0];
	reg [82:0] body_die [73:0];
	reg [82:0] feet_normal [13:0];
	reg [82:0] feet_left [13:0];
	reg [82:0] feet_right [13:0];
	
	reg [82:0] body [73:0];
	reg [82:0] feet [13:0];
	
	initial begin
		body_normal[0] = 82'b0000000000_0000000000_0000000000_0000000000_0000000011_1111111111_1111111111_1111111100_00;
        body_normal[1] = 82'b0000000000_0000000000_0000000000_0000000000_0000000011_1111111111_1111111111_1111111100_00;
        body_normal[2] = 82'b0000000000_0000000000_0000000000_0000000000_0000000011_1111111111_1111111111_1111111100_00;
        body_normal[3] = 82'b0000000000_0000000000_0000000000_0000000000_0000000011_1111111111_1111111111_1111111100_00;
        body_normal[4] = 82'b0000000000_0000000000_0000000000_0000000000_0000111111_1111111111_1111111111_1111111111_11;
        body_normal[5] = 82'b0000000000_0000000000_0000000000_0000000000_0000111111_1111111111_1111111111_1111111111_11;
        body_normal[6] = 82'b0000000000_0000000000_0000000000_0000000000_0000111111_1111111111_1111111111_1111111111_11;
        body_normal[7] = 82'b0000000000_0000000000_0000000000_0000000000_0000111111_1111111111_1111111111_1111111111_11;
        body_normal[8] = 82'b0000000000_0000000000_0000000000_0000000000_0000111111_1100011111_1111111111_1111111111_11;
        body_normal[9] = 82'b0000000000_0000000000_0000000000_0000000000_0000111111_1100011111_1111111111_1111111111_11;
        body_normal[10] = 82'b0000000000_0000000000_0000000000_0000000000_0000111111_1100011111_1111111111_1111111111_11;
        body_normal[11] = 82'b0000000000_0000000000_0000000000_0000000000_0000111111_1111111111_1111111111_1111111111_11;
        body_normal[12] = 82'b0000000000_0000000000_0000000000_0000000000_0000111111_1111111111_1111111111_1111111111_11;
        body_normal[13] = 82'b0000000000_0000000000_0000000000_0000000000_0000111111_1111111111_1111111111_1111111111_11;
        body_normal[14] = 82'b0000000000_0000000000_0000000000_0000000000_0000111111_1111111111_1111111111_1111111111_11;
        body_normal[15] = 82'b0000000000_0000000000_0000000000_0000000000_0000111111_1111111111_1111111111_1111111111_11;
        body_normal[16] = 82'b0000000000_0000000000_0000000000_0000000000_0000111111_1111111111_1111111111_1111111111_11;
        body_normal[17] = 82'b0000000000_0000000000_0000000000_0000000000_0000111111_1111111111_1111111111_1111111111_11;
        body_normal[18] = 82'b0000000000_0000000000_0000000000_0000000000_0000111111_1111111111_1111111111_1111111111_11;
        body_normal[19] = 82'b0000000000_0000000000_0000000000_0000000000_0000111111_1111111111_1111111111_1111111111_11;
        body_normal[20] = 82'b0000000000_0000000000_0000000000_0000000000_0000111111_1111111111_1111111111_1111111111_11;
        body_normal[21] = 82'b0000000000_0000000000_0000000000_0000000000_0000111111_1111111111_1111111111_1111111111_11;
        body_normal[22] = 82'b0000000000_0000000000_0000000000_0000000000_0000111111_1111111111_1111111111_1111111111_11;
        body_normal[23] = 82'b0000000000_0000000000_0000000000_0000000000_0000111111_1111111111_1110000000_0000000000_00;
        body_normal[24] = 82'b0000000000_0000000000_0000000000_0000000000_0000111111_1111111111_1110000000_0000000000_00;
        body_normal[25] = 82'b0000000000_0000000000_0000000000_0000000000_0000111111_1111111111_1110000000_0000000000_00;
        body_normal[26] = 82'b1111000000_0000000000_0000000000_0000000000_1111111111_1111111111_1111111111_1111111100_00;
        body_normal[27] = 82'b1111000000_0000000000_0000000000_0000000000_1111111111_1111111111_1111111111_1111111100_00;
        body_normal[28] = 82'b1111000000_0000000000_0000000000_0000001111_1111111111_1111110000_0000000000_0000000000_00;
        body_normal[29] = 82'b1111000000_0000000000_0000000000_0000001111_1111111111_1111110000_0000000000_0000000000_00;
        body_normal[30] = 82'b1111000000_0000000000_0000000000_0000111111_1111111111_1111110000_0000000000_0000000000_00;
        body_normal[31] = 82'b1111000000_0000000000_0000000000_0000111111_1111111111_1111110000_0000000000_0000000000_00;
        body_normal[32] = 82'b1111110000_0000000000_0000000000_0011111111_1111111111_1111110000_0000000000_0000000000_00;
        body_normal[33] = 82'b1111110000_0000000000_0000000000_0011111111_1111111111_1111110000_0000000000_0000000000_00;
        body_normal[34] = 82'b1111111100_0000000000_0000000000_1111111111_1111111111_1111110000_0000000000_0000000000_00;
        body_normal[35] = 82'b1111111100_0000000000_0000000000_1111111111_1111111111_1111110000_0000000000_0000000000_00;
        body_normal[36] = 82'b1111111111_0000000000_0000001111_1111111111_1111111111_1111110000_0000000000_0000000000_00;
        body_normal[37] = 82'b1111111111_0000000000_0000001111_1111111111_1111111111_1111110000_0000000000_0000000000_00;
        body_normal[38] = 82'b1111111111_1100000000_0000111111_1111111111_1111111111_1111111111_1111000000_0000000000_00;
        body_normal[39] = 82'b1111111111_1100000000_0000111111_1111111111_1111111111_1111111111_1111000000_0000000000_00;
        body_normal[40] = 82'b1111111111_1111000000_1111111111_1111111111_1111111111_1111111111_1111000000_0000000000_00;
        body_normal[41] = 82'b1111111111_1111000000_1111111111_1111111111_1111111111_1111111111_1111000000_0000000000_00;
        body_normal[42] = 82'b1111111111_1111111111_1111111111_1111111111_1111111111_1111110000_1111000000_0000000000_00;
        body_normal[43] = 82'b1111111111_1111111111_1111111111_1111111111_1111111111_1111110000_1111000000_0000000000_00;
        body_normal[44] = 82'b1111111111_1111111111_1111111111_1111111111_1111111111_1111110000_1111000000_0000000000_00;
        body_normal[45] = 82'b1111111111_1111111111_1111111111_1111111111_1111111111_1111110000_1111000000_0000000000_00;
        body_normal[46] = 82'b1111111111_1111111111_1111111111_1111111111_1111111111_1111110000_0000000000_0000000000_00;
        body_normal[47] = 82'b1111111111_1111111111_1111111111_1111111111_1111111111_1111110000_0000000000_0000000000_00;
        body_normal[48] = 82'b1111111111_1111111111_1111111111_1111111111_1111111111_1111110000_0000000000_0000000000_00;
        body_normal[49] = 82'b1111111111_1111111111_1111111111_1111111111_1111111111_1111110000_0000000000_0000000000_00;
        body_normal[50] = 82'b1111111111_1111111111_1111111111_1111111111_1111111111_1111110000_0000000000_0000000000_00;
        body_normal[51] = 82'b1111111111_1111111111_1111111111_1111111111_1111111111_1111110000_0000000000_0000000000_00;
        body_normal[52] = 82'b1111111111_1111111111_1111111111_1111111111_1111111111_1111110000_0000000000_0000000000_00;
        body_normal[53] = 82'b1111111111_1111111111_1111111111_1111111111_1111111111_1111110000_0000000000_0000000000_00;
        body_normal[54] = 82'b0011111111_1111111111_1111111111_1111111111_1111111111_1111110000_0000000000_0000000000_00;
        body_normal[55] = 82'b0011111111_1111111111_1111111111_1111111111_1111111111_1111110000_0000000000_0000000000_00;
        body_normal[56] = 82'b0000111111_1111111111_1111111111_1111111111_1111111111_1111110000_0000000000_0000000000_00;
        body_normal[57] = 82'b0000111111_1111111111_1111111111_1111111111_1111111111_1111110000_0000000000_0000000000_00;
        body_normal[58] = 82'b0000001111_1111111111_1111111111_1111111111_1111111111_1111110000_0000000000_0000000000_00;
        body_normal[59] = 82'b0000001111_1111111111_1111111111_1111111111_1111111111_1111110000_0000000000_0000000000_00;
        body_normal[60] = 82'b0000000011_1111111111_1111111111_1111111111_1111111111_1111110000_0000000000_0000000000_00;
        body_normal[61] = 82'b0000000011_1111111111_1111111111_1111111111_1111111111_1111110000_0000000000_0000000000_00;
        body_normal[62] = 82'b0000000000_1111111111_1111111111_1111111111_1111111111_1111000000_0000000000_0000000000_00;
        body_normal[63] = 82'b0000000000_1111111111_1111111111_1111111111_1111111111_1111000000_0000000000_0000000000_00;
        body_normal[64] = 82'b0000000000_0011111111_1111111111_1111111111_1111111111_1100000000_0000000000_0000000000_00;
        body_normal[65] = 82'b0000000000_0011111111_1111111111_1111111111_1111111111_1100000000_0000000000_0000000000_00;
        body_normal[66] = 82'b0000000000_0000111111_1111111111_1111111111_1111111111_0000000000_0000000000_0000000000_00;
        body_normal[67] = 82'b0000000000_0000111111_1111111111_1111111111_1111111111_0000000000_0000000000_0000000000_00;
        body_normal[68] = 82'b0000000000_0000001111_1111111111_1111111111_1111111100_0000000000_0000000000_0000000000_00;
        body_normal[69] = 82'b0000000000_0000001111_1111111111_1111111111_1111111100_0000000000_0000000000_0000000000_00;
        body_normal[70] = 82'b0000000000_0000000011_1111111111_1111111111_1111110000_0000000000_0000000000_0000000000_00;
        body_normal[71] = 82'b0000000000_0000000011_1111111111_1111111111_1111110000_0000000000_0000000000_0000000000_00;
        body_normal[72] = 82'b0000000000_0000000000_1111111111_1111111111_1111000000_0000000000_0000000000_0000000000_00;
        body_normal[73] = 82'b0000000000_0000000000_1111111111_1111111111_1111000000_0000000000_0000000000_0000000000_00;
		
		body_die[0] = 82'b0000000000_0000000000_0000000000_0000000000_0000000011_1111111111_1111111111_1111111100_00;
        body_die[1] = 82'b0000000000_0000000000_0000000000_0000000000_0000000011_1111111111_1111111111_1111111100_00;
        body_die[2] = 82'b0000000000_0000000000_0000000000_0000000000_0000000011_1111111111_1111111111_1111111100_00;
        body_die[3] = 82'b0000000000_0000000000_0000000000_0000000000_0000000011_1111111111_1111111111_1111111100_00;
        body_die[4] = 82'b0000000000_0000000000_0000000000_0000000000_0000111111_1111111111_1111111111_1111111111_11;
        body_die[5] = 82'b0000000000_0000000000_0000000000_0000000000_0000111111_1111111111_1111111111_1111111111_11;
        body_die[6] = 82'b0000000000_0000000000_0000000000_0000000000_0000111111_0000001111_1111111111_1111111111_11;
        body_die[7] = 82'b0000000000_0000000000_0000000000_0000000000_0000111111_0000001111_1111111111_1111111111_11;
        body_die[8] = 82'b0000000000_0000000000_0000000000_0000000000_0000111111_0011001111_1111111111_1111111111_11;
        body_die[9] = 82'b0000000000_0000000000_0000000000_0000000000_0000111111_0011001111_1111111111_1111111111_11;
        body_die[10] = 82'b0000000000_0000000000_0000000000_0000000000_0000111111_0000001111_1111111111_1111111111_11;
        body_die[11] = 82'b0000000000_0000000000_0000000000_0000000000_0000111111_0000001111_1111111111_1111111111_11;
        body_die[12] = 82'b0000000000_0000000000_0000000000_0000000000_0000111111_1111111111_1111111111_1111111111_11;
        body_die[13] = 82'b0000000000_0000000000_0000000000_0000000000_0000111111_1111111111_1111111111_1111111111_11;
        body_die[14] = 82'b0000000000_0000000000_0000000000_0000000000_0000111111_1111111111_1111111111_1111111111_11;
        body_die[15] = 82'b0000000000_0000000000_0000000000_0000000000_0000111111_1111111111_1111111111_1111111111_11;
        body_die[16] = 82'b0000000000_0000000000_0000000000_0000000000_0000111111_1111111111_1111111111_1111111111_11;
        body_die[17] = 82'b0000000000_0000000000_0000000000_0000000000_0000111111_1111111111_1111111111_1111111111_11;
        body_die[18] = 82'b0000000000_0000000000_0000000000_0000000000_0000111111_1111111111_1111111111_1111111111_11;
        body_die[19] = 82'b0000000000_0000000000_0000000000_0000000000_0000111111_1111111111_1111111111_1111111111_11;
        body_die[20] = 82'b0000000000_0000000000_0000000000_0000000000_0000111111_1111111111_1111111111_1111111111_11;
        body_die[21] = 82'b0000000000_0000000000_0000000000_0000000000_0000111111_1111111111_1111111111_1111111111_11;
        body_die[22] = 82'b0000000000_0000000000_0000000000_0000000000_0000111111_1111111111_1111111111_1111111111_11;
        body_die[23] = 82'b0000000000_0000000000_0000000000_0000000000_0000111111_1111111111_1111111111_1111111111_11;
        body_die[24] = 82'b0000000000_0000000000_0000000000_0000000000_0000111111_1111111111_1111111111_1111111100_00;
        body_die[25] = 82'b0000000000_0000000000_0000000000_0000000000_0000111111_1111111111_1111111111_1111111100_00;
        body_die[26] = 82'b1111000000_0000000000_0000000000_0000000000_1111111111_1111111111_1111111111_1111111100_00;
        body_die[27] = 82'b1111000000_0000000000_0000000000_0000000000_1111111111_1111111111_1111111111_1111111100_00;
        body_die[28] = 82'b1111000000_0000000000_0000000000_0000001111_1111111111_1111110000_0000000000_0000000000_00;
        body_die[29] = 82'b1111000000_0000000000_0000000000_0000001111_1111111111_1111110000_0000000000_0000000000_00;
        body_die[30] = 82'b1111000000_0000000000_0000000000_0000111111_1111111111_1111110000_0000000000_0000000000_00;
        body_die[31] = 82'b1111000000_0000000000_0000000000_0000111111_1111111111_1111110000_0000000000_0000000000_00;
        body_die[32] = 82'b1111110000_0000000000_0000000000_0011111111_1111111111_1111110000_0000000000_0000000000_00;
        body_die[33] = 82'b1111110000_0000000000_0000000000_0011111111_1111111111_1111110000_0000000000_0000000000_00;
        body_die[34] = 82'b1111111100_0000000000_0000000000_1111111111_1111111111_1111110000_0000000000_0000000000_00;
        body_die[35] = 82'b1111111100_0000000000_0000000000_1111111111_1111111111_1111110000_0000000000_0000000000_00;
        body_die[36] = 82'b1111111111_0000000000_0000001111_1111111111_1111111111_1111110000_0000000000_0000000000_00;
        body_die[37] = 82'b1111111111_0000000000_0000001111_1111111111_1111111111_1111110000_0000000000_0000000000_00;
        body_die[38] = 82'b1111111111_1100000000_0000111111_1111111111_1111111111_1111111111_1111000000_0000000000_00;
        body_die[39] = 82'b1111111111_1100000000_0000111111_1111111111_1111111111_1111111111_1111000000_0000000000_00;
        body_die[40] = 82'b1111111111_1111000000_1111111111_1111111111_1111111111_1111111111_1111000000_0000000000_00;
        body_die[41] = 82'b1111111111_1111000000_1111111111_1111111111_1111111111_1111111111_1111000000_0000000000_00;
        body_die[42] = 82'b1111111111_1111111111_1111111111_1111111111_1111111111_1111110000_1111000000_0000000000_00;
        body_die[43] = 82'b1111111111_1111111111_1111111111_1111111111_1111111111_1111110000_1111000000_0000000000_00;
        body_die[44] = 82'b1111111111_1111111111_1111111111_1111111111_1111111111_1111110000_1111000000_0000000000_00;
        body_die[45] = 82'b1111111111_1111111111_1111111111_1111111111_1111111111_1111110000_1111000000_0000000000_00;
        body_die[46] = 82'b1111111111_1111111111_1111111111_1111111111_1111111111_1111110000_0000000000_0000000000_00;
        body_die[47] = 82'b1111111111_1111111111_1111111111_1111111111_1111111111_1111110000_0000000000_0000000000_00;
        body_die[48] = 82'b1111111111_1111111111_1111111111_1111111111_1111111111_1111110000_0000000000_0000000000_00;
        body_die[49] = 82'b1111111111_1111111111_1111111111_1111111111_1111111111_1111110000_0000000000_0000000000_00;
        body_die[50] = 82'b1111111111_1111111111_1111111111_1111111111_1111111111_1111110000_0000000000_0000000000_00;
        body_die[51] = 82'b1111111111_1111111111_1111111111_1111111111_1111111111_1111110000_0000000000_0000000000_00;
        body_die[52] = 82'b1111111111_1111111111_1111111111_1111111111_1111111111_1111110000_0000000000_0000000000_00;
        body_die[53] = 82'b1111111111_1111111111_1111111111_1111111111_1111111111_1111110000_0000000000_0000000000_00;
        body_die[54] = 82'b0011111111_1111111111_1111111111_1111111111_1111111111_1111110000_0000000000_0000000000_00;
        body_die[55] = 82'b0011111111_1111111111_1111111111_1111111111_1111111111_1111110000_0000000000_0000000000_00;
        body_die[56] = 82'b0000111111_1111111111_1111111111_1111111111_1111111111_1111110000_0000000000_0000000000_00;
        body_die[57] = 82'b0000111111_1111111111_1111111111_1111111111_1111111111_1111110000_0000000000_0000000000_00;
        body_die[58] = 82'b0000001111_1111111111_1111111111_1111111111_1111111111_1111110000_0000000000_0000000000_00;
        body_die[59] = 82'b0000001111_1111111111_1111111111_1111111111_1111111111_1111110000_0000000000_0000000000_00;
        body_die[60] = 82'b0000000011_1111111111_1111111111_1111111111_1111111111_1111110000_0000000000_0000000000_00;
        body_die[61] = 82'b0000000011_1111111111_1111111111_1111111111_1111111111_1111110000_0000000000_0000000000_00;
        body_die[62] = 82'b0000000000_1111111111_1111111111_1111111111_1111111111_1111000000_0000000000_0000000000_00;
        body_die[63] = 82'b0000000000_1111111111_1111111111_1111111111_1111111111_1111000000_0000000000_0000000000_00;
        body_die[64] = 82'b0000000000_0011111111_1111111111_1111111111_1111111111_1100000000_0000000000_0000000000_00;
        body_die[65] = 82'b0000000000_0011111111_1111111111_1111111111_1111111111_1100000000_0000000000_0000000000_00;
        body_die[66] = 82'b0000000000_0000111111_1111111111_1111111111_1111111111_0000000000_0000000000_0000000000_00;
        body_die[67] = 82'b0000000000_0000111111_1111111111_1111111111_1111111111_0000000000_0000000000_0000000000_00;
        body_die[68] = 82'b0000000000_0000001111_1111111111_1111111111_1111111100_0000000000_0000000000_0000000000_00;
        body_die[69] = 82'b0000000000_0000001111_1111111111_1111111111_1111111100_0000000000_0000000000_0000000000_00;
        body_die[70] = 82'b0000000000_0000000011_1111111111_1111111111_1111110000_0000000000_0000000000_0000000000_00;
        body_die[71] = 82'b0000000000_0000000011_1111111111_1111111111_1111110000_0000000000_0000000000_0000000000_00;
        body_die[72] = 82'b0000000000_0000000000_1111111111_1111111111_1111000000_0000000000_0000000000_0000000000_00;
        body_die[73] = 82'b0000000000_0000000000_1111111111_1111111111_1111000000_0000000000_0000000000_0000000000_00;
		
		feet_normal[0] = 82'b0000000000_0000000000_1111111111_1100001111_1111000000_0000000000_0000000000_0000000000_00;
        feet_normal[1] = 82'b0000000000_0000000000_1111111111_1100001111_1111000000_0000000000_0000000000_0000000000_00;
        feet_normal[2] = 82'b0000000000_0000000000_1111111100_0000000000_1111000000_0000000000_0000000000_0000000000_00;
        feet_normal[3] = 82'b0000000000_0000000000_1111111100_0000000000_1111000000_0000000000_0000000000_0000000000_00;
        feet_normal[4] = 82'b0000000000_0000000000_1111111100_0000000000_1111000000_0000000000_0000000000_0000000000_00;
        feet_normal[5] = 82'b0000000000_0000000000_1111110000_0000000000_1111000000_0000000000_0000000000_0000000000_00;
        feet_normal[6] = 82'b0000000000_0000000000_1111000000_0000000000_1111000000_0000000000_0000000000_0000000000_00;
        feet_normal[7] = 82'b0000000000_0000000000_1111000000_0000000000_1111000000_0000000000_0000000000_0000000000_00;
        feet_normal[8] = 82'b0000000000_0000000000_1111000000_0000000000_1111000000_0000000000_0000000000_0000000000_00;
        feet_normal[9] = 82'b0000000000_0000000000_1111000000_0000000000_1111000000_0000000000_0000000000_0000000000_00;
        feet_normal[10] = 82'b0000000000_0000000000_1111111100_0000000000_1111111100_0000000000_0000000000_0000000000_00;
        feet_normal[11] = 82'b0000000000_0000000000_1111111100_0000000000_1111111100_0000000000_0000000000_0000000000_00;
        feet_normal[12] = 82'b0000000000_0000000000_1111111100_0000000000_1111111100_0000000000_0000000000_0000000000_00;
        feet_normal[13] = 82'b0000000000_0000000000_1111111100_0000000000_1111111100_0000000000_0000000000_0000000000_00;
		
		feet_left[0] = 82'b0000000000_0000000000_1111111100_0000001111_1111000000_0000000000_0000000000_0000000000_00;
		feet_left[1] = 82'b0000000000_0000000000_1111111100_0000001111_1111000000_0000000000_0000000000_0000000000_00;
		feet_left[2] = 82'b0000000000_0000000000_1111111100_0000000000_1111000000_0000000000_0000000000_0000000000_00;
		feet_left[3] = 82'b0000000000_0000000000_0011111111_1111000000_1111000000_0000000000_0000000000_0000000000_00;
		feet_left[4] = 82'b0000000000_0000000000_0011111111_1111000000_1111000000_0000000000_0000000000_0000000000_00;
		feet_left[5] = 82'b0000000000_0000000000_0000000000_0000000000_1111000000_0000000000_0000000000_0000000000_00;
		feet_left[6] = 82'b0000000000_0000000000_0000000000_0000000000_1111000000_0000000000_0000000000_0000000000_00;
		feet_left[7] = 82'b0000000000_0000000000_0000000000_0000000000_1111000000_0000000000_0000000000_0000000000_00;
		feet_left[8] = 82'b0000000000_0000000000_0000000000_0000000000_1111000000_0000000000_0000000000_0000000000_00;
		feet_left[9] = 82'b0000000000_0000000000_0000000000_0000000000_1111000000_0000000000_0000000000_0000000000_00;
		feet_left[10] = 82'b0000000000_0000000000_0000000000_0000000000_1111111100_0000000000_0000000000_0000000000_00;
		feet_left[11] = 82'b0000000000_0000000000_0000000000_0000000000_1111111100_0000000000_0000000000_0000000000_00;
		feet_left[12] = 82'b0000000000_0000000000_0000000000_0000000000_1111111100_0000000000_0000000000_0000000000_00;
		feet_left[13] = 82'b0000000000_0000000000_0000000000_0000000000_1111111100_0000000000_0000000000_0000000000_00;
		
		feet_right[0] = 82'b0000000000_0000000000_1111111111_1100000000_1111000000_0000000000_0000000000_0000000000_00;
        feet_right[1] = 82'b0000000000_0000000000_1111111111_1100000000_1111000000_0000000000_0000000000_0000000000_00;
        feet_right[2] = 82'b0000000000_0000000000_1111111100_0000000000_1111111111_0000000000_0000000000_0000000000_00;
        feet_right[3] = 82'b0000000000_0000000000_1111111100_0000000000_1111111111_0000000000_0000000000_0000000000_00;
        feet_right[4] = 82'b0000000000_0000000000_1111111100_0000000000_0000000000_0000000000_0000000000_0000000000_00;
        feet_right[5] = 82'b0000000000_0000000000_1111110000_0000000000_0000000000_0000000000_0000000000_0000000000_00;
        feet_right[6] = 82'b0000000000_0000000000_1111000000_0000000000_0000000000_0000000000_0000000000_0000000000_00;
        feet_right[7] = 82'b0000000000_0000000000_1111000000_0000000000_0000000000_0000000000_0000000000_0000000000_00;
        feet_right[8] = 82'b0000000000_0000000000_1111000000_0000000000_0000000000_0000000000_0000000000_0000000000_00;
        feet_right[9] = 82'b0000000000_0000000000_1111000000_0000000000_0000000000_0000000000_0000000000_0000000000_00;
        feet_right[10] = 82'b0000000000_0000000000_1111111100_0000000000_0000000000_0000000000_0000000000_0000000000_00;
        feet_right[11] = 82'b0000000000_0000000000_1111111100_0000000000_0000000000_0000000000_0000000000_0000000000_00;
        feet_right[12] = 82'b0000000000_0000000000_1111111100_0000000000_0000000000_0000000000_0000000000_0000000000_00;
        feet_right[13] = 82'b0000000000_0000000000_1111111100_0000000000_0000000000_0000000000_0000000000_0000000000_00;
	end
/* --------------------------------------------------------------------------------------------------------------------------- */
	
	// === 實例化偵測按鈕的module(改成在top module實例) ===
	/*
	wire key_flag;
	wire key_value;
	key_debounce u_key_debounce(
		.clk(lcd_pclk), 
		.rst_n(rst_n), 
		.key(key),
		.key_flag(key_flag), 
		.key_value(key_value)
	);*/
	
/* --------------------------------------------------------------------------------------------------------------------------- */

	// === 決定輸入的pixel 是否要印出恐龍的黑色 ===
	parameter DINO_X = 20;
	parameter DINO_Y = 360;
    parameter BODY_H = 74;
    parameter FEET_H = 14;
    parameter DINO_H = BODY_H + FEET_H;  // 總高 88
	parameter DINO_W = 83;
	reg [9:0] jump_height;
	
	// === 相對 pixel 位置 ===
    wire [6:0] rel_x = pixel_xpos - DINO_X;
    wire [6:0] rel_y = pixel_ypos - (DINO_Y - jump_height);

	wire in_range = (pixel_xpos >= DINO_X) && (pixel_xpos < DINO_X + DINO_W) &&
                    (pixel_ypos >= (DINO_Y - jump_height)) && (pixel_ypos < (DINO_Y - jump_height) + DINO_H);

    // === bitmap 查表邏輯 ===
    wire body_bit = (rel_y < BODY_H) ? body[rel_y][82 - rel_x] : 1'b0;
    wire feet_bit = (rel_y >= BODY_H && rel_y < DINO_H) ? feet[rel_y - BODY_H][82 - rel_x] : 1'b0;
	
	assign dino_draw = in_range && (body_bit || feet_bit);
	
	
	integer i;
	always @(*) begin
		for (i = 0; i < 74; i = i + 1) begin
			case (dino_state)
				normal: begin
					body[i] = body_normal[i];
				end
				jump: begin
					body[i] = body_normal[i];
				end
				run_left: begin
					body[i] = body_normal[i];
				end
				run_right: begin
					body[i] = body_normal[i];
				end
				die: begin
					body[i] = body_die[i];
				end
				default: begin
					body[i] = body_normal[i];
				end
			endcase
		end
		
		for (i = 0; i < 14; i = i + 1) begin
			case (dino_state)
				normal: begin
					feet[i] = feet_normal[i];
				end
				jump: begin
					feet[i] = feet_normal[i];
				end
				run_left: begin
					feet[i] = feet_left[i];
				end
				run_right: begin
					feet[i] = feet_right[i];
				end
				die: begin
					feet[i] = feet_normal[i];
				end
				default: begin
					feet[i] = feet_normal[i];
				end
			endcase
		end
	end
	
/* --------------------------------------------------------------------------------------------------------------------------- */

	// === 更新恐龍狀態和位置(跳躍 奔跑 掛掉) ===
	parameter normal = 3'd0;
	parameter run_left = 3'd1;
	parameter run_right = 3'd2;
	parameter jump = 3'd3;
	parameter die = 3'd4;
	reg [2:0] dino_state;
	reg [7:0] jump_time;
	parameter JUMP_TIME_LIMIT = 8'd56;

	// === 100HZ時鐘 用於更新跳躍位置 ===
	reg [17:0] clk_100_counter;
	parameter clk_100_CNT = 18'd125000;
	
	always @(posedge lcd_pclk or negedge rst_n) begin
		if(!rst_n) begin
			clk_100 <= 1'b0;
			clk_100_counter <= 18'd0;
		end
		else begin
			if(clk_100_counter < clk_100_CNT - 1'b1) 
				clk_100_counter <= clk_100_counter + 1'b1;
			else begin
				clk_100_counter <= 18'd0;
				clk_100 <= ~clk_100;
			end
		end
	end
	
	// === 10HZ時鐘 用於更新左右腳跑步 ===
	reg clk_10;
	reg clk_10_prev;
	reg [3:0] clk_10_counter;
	parameter clk_10_CNT = 4'd5;
	
	always @(posedge clk_100 or negedge rst_n) begin
		if(!rst_n) begin
			clk_10 <= 1'b0;
			clk_10_counter <= 4'd0;
		end
		else begin
			if(clk_10_counter < clk_10_CNT - 1'b1) 
				clk_10_counter <= clk_10_counter + 1'b1;
			else begin
				clk_10_counter <= 4'd0;
				clk_10 <= ~clk_10;
			end
		end
	end
	
	// === 更新恐龍state以及圖案長相 ===
	always @(posedge lcd_pclk or negedge rst_n) begin
		if(!rst_n) begin
			dino_state <= normal;
			clk_10_prev <= 1'b0;
		end
		else if(is_dying) begin
			dino_state <= die;
		end
		else begin
			// 更新 clk_10_prev
			clk_10_prev <= clk_10;

			if(dino_state == jump) begin
				if(jump_time >= JUMP_TIME_LIMIT - 1)
					dino_state <= run_left;
				else
					dino_state <= jump;
			end
			else if(key_flag && (~key_value)) begin
				dino_state <= jump;
			end
			else if(clk_10 && ~clk_10_prev) begin
				case(dino_state)
					normal:    dino_state <= normal;
					run_left:  dino_state <= run_right;
					run_right: dino_state <= run_left;
					default:   dino_state <= dino_state;
				endcase
			end
			else begin
				dino_state <= dino_state;
			end
		end
	end

	// === 即時更新恐龍高度 不是jump狀態下會是0 (會用基準點 - 高度) === 
	always @(*) begin
		/*if (((jump_time * 15) - (jump_time * jump_time) / 2) > 0)
			jump_height = (jump_time * 15) - (jump_time * jump_time) / 2;
		else
			jump_height = 0;*/
		jump_height = (jump_time * 14) - (jump_time * jump_time) / 4;
	end

	// === jump狀態下的持續滯空時間 === 
	always @(posedge clk_100 or negedge rst_n) begin
		if (!rst_n)
			jump_time <= 0;
		else if(is_living) begin
			if (dino_state == jump)
				jump_time <= jump_time + 1;
			else
				jump_time <= 0;
		end
	end
/* --------------------------------------------------------------------------------------------------------------------------- */
	
endmodule