module ground(
    input	lcd_pclk,
	input	clk_100,
    input	rst_n,
    input	[10:0]  pixel_xpos,
    input	[10:0]  pixel_ypos,
	input	is_living,
	input	[3:0] move_rate,

    output reg ground_draw
);

	reg [159:0] ground [9:0];
	initial begin
		ground[0]<=160'b0000000000_0000000000_0000000000_0000000000_1111100000_0000000000_0000000000_1111111111_0000000000_0000000000_0000000000_1111111111_0000000000_0000000000_0000000000_1111111111;
		ground[1]<=160'b1111100000_1111111111_1111111111_1111111111_1111111111_1111111111_1111111111_0000000000_1111111111_1111111111_1111111111_0000000000_1111111111_1111111111_1111111111_0000000000;
		ground[2]<=160'b0000011111_0000000000_0000000000_0000000000_0000000000_1111000000_0000000000_0000000000_0000000000_0000000000_0001111110_0000000000_0000000000_0000000000_0000000000_0000000000;
        ground[3]<=160'b0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000;
        ground[4]<=160'b0000000000_0111000000_0000000000_0000000011_1000000000_0000000000_0000000000_0000000000_0000000110_0000000000_0000000000_0111000000_0000000000_0000000000_0000000000_0000000000;
        ground[5]<=160'b0000000000_0000000000_0000000000_0000000000_0000110000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000111000_0000000000_0000000000_0000000000;
        ground[6]<=160'b0000000000_0100000000_0000000000_0000110000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0011000000;
        ground[7]<=160'b0000000000_0000000000_0000011100_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0011110000_0000000000_0000000000_0000000000_0000000000_0000000000;
        ground[8]<=160'b0000000010_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0011000000_0000000000_0000000000_0000000000_0000000000_0000000000_1110000000_0000000000_0000000000;
        ground[9]<=160'b0000000000_0111000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000001000;
	end
	
	// === 地板參數 ===
    parameter GND_X = 0;         // 地板起始 X
    parameter GND_Y = 435;       // 地板起始 Y
    parameter GND_W = 800;       // 實際畫滿 800 pixels
    parameter GND_H = 10;

    // === 顯示控制邏輯(靜態) ===
    /*
	always @(*) begin
        if (pixel_xpos >= GND_X && pixel_xpos < GND_X + GND_W &&
            pixel_ypos >= GND_Y && pixel_ypos < GND_Y + GND_H) begin

            // X 座標超過 160，就取餘數，達到重複 pattern 效果
            ground_draw = ground[pixel_ypos - GND_Y][(pixel_xpos - GND_X) % 160];
        end 
		else begin
            ground_draw = 1'b0;
        end
    end		*/
	
	reg [7:0] scroll_offset;
	always @(posedge clk_100 or negedge rst_n) begin
		if(!rst_n)
			scroll_offset <= 8'd0;
		else if(is_living)
			scroll_offset <= (scroll_offset + move_rate) % 8'd160;
	end
	
	always @(*) begin
        if (pixel_xpos >= GND_X && pixel_xpos < GND_X + GND_W &&
            pixel_ypos >= GND_Y && pixel_ypos < GND_Y + GND_H) begin

            // X 座標超過 160，就取餘數，達到重複 pattern 效果
            ground_draw = ground[pixel_ypos - GND_Y][(pixel_xpos + scroll_offset - GND_X) % 160];
        end 
		else begin
            ground_draw = 1'b0;
        end
    end	

endmodule